//+++++++++++++++++++++++=++++++++++++++++++++++++++
//Author:			
//
//--------- ----------------------------------------
//+Verison+  								Describe
//--------- ----------------------------------------
//   0.0								Initial Verison
//--------- ----------------------------------------
//+++++++++++++++++++++++=++++++++++++++++++++++++++
									

module tb_top;




initial begin
	$fsdbDumpfile("tb_top.fsdb");
	$fsdbDumpvars();
end

endmodule
